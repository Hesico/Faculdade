module ou(
			input [3:0] A,B,
			output[3:0] ouAB
			);
			
or or0(ouAB[0], A[0],B[0]);
or or1(ouAB[1], A[1],B[1]);
or or2(ouAB[2], A[2],B[2]);
or or3(ouAB[3], A[3],B[3]);			
			  
endmodule 